`timescale 1ns / 1ps

module AND_GATE(output Y, input A,B); //Declaring AND Gate Module with Y as OUTPUT and A,B as INPUT.

and F1(Y,A,B);                        //Using inbuilt 'and' gate.

endmodule
