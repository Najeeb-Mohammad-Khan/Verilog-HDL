`timescale 1ns / 1ps

module NOT_GATE(output Y,input A);   ////Declaring NOT Gate Module with Y as OUTPUT and A as INPUT.

not F1(Y,A);   // Using inbuilt 'not' gate.

endmodule
