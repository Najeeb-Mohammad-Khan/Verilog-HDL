`timescale 1ns / 1ps

module OR_GATE(output Y, input A,B);		//Declaring OR_GATE module with Y as OUTPUT and A,B as INPUT.

or F1(Y,A,B);		//Using inbuilt 'OR' Gate.

endmodule
